//`define SIMULATION

`define SOFTMC_STREAM_WIDTH 256
`define SOFTMC_STREAM_KEEP  32

`define DQ_WIDTH        64
`define ODT_WIDTH       1
`define CS_WIDTH        1
`define CKE_WIDTH       1
`define CK_WIDTH        1
`define ROW_ADDR_WIDTH  14

`define BANK_WIDTH      3
`define ROW_WIDTH       16