// `define ENABLE_DLL_TOGGLER
`define DQ_WIDTH 64
// DIMM related
`define ODT_WIDTH  1
`define CS_WIDTH   1
`define CKE_WIDTH  1
`define CK_WIDTH   1